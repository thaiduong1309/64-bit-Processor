module CPU();
	logic [63:0]WriteData;
	logic [4:0]ReadRegister1, ReadRegister2, WriteRegister;
	logic clk,RegWrite,reset;
	logic [63:0]ReadData1, ReadData2;
	logic		[2:0]		cntrl;
	logic	[63:0]	result;
	logic	negative, zero, overflow, carry_out;
	logic		[31:0]	instruction




endmodule