library verilog;
use verilog.vl_types.all;
entity DFF_REG_testbench is
end DFF_REG_testbench;
